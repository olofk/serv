localparam [1:0]
  CSR_MSCRATCH = 2'b00,
  CSR_MTVEC    = 2'b01,
  CSR_MEPC     = 2'b10,
  CSR_MTVAL    = 2'b11;
